`timescale 1ns/10ps
`include "./median.v"
module tb;

reg    [7:0] a0, a1, a2;
wire   [7:0] out;

median m0 (a0, a1, a2, out);

initial begin
    a0=8'b00000000 ;a1=8'b00000000 ;a2=8'b00000000;
#10	a0=8'b10000000 ;a1=8'b00010000 ;a2=8'b00000001; //case 3'b000
#60 a0=8'b00100000 ;a1=8'b01000000 ;a2=8'b00000100; //case 3'b001
#110 a0=8'b00000010 ;a1=8'b00100000 ;a2=8'b00001000; //cade 3'b011  
#150 a0=8'b01000000 ;a1=8'b00001000 ;a2=8'b00010000; //case 3'b100
#210 a0=8'b00001000 ;a1=8'b00000010 ;a2=8'b01000000; //case 3'b110
#260 a0=8'b00000001 ;a1=8'b00001000 ;a2=8'b10000000; //case 3'b111
#310 a0=8'b00000100 ;a1=8'b00000100 ;a2=8'b00100000; //a0=a1
#360 a0=8'b00100000 ;a1=8'b00010000 ;a2=8'b00010000; //a1=a2
#410 a0=8'b10000000 ;a2=8'b00000001 ;a2=8'b10000000; //a0=a2
#460 a0=8'b00000000 ;a2=8'b00000001 ;a2=8'b10000000; //a0=b'd0
#510 a0=8'b10000000 ;a1=8'b00000000 ;a2=8'b00000001; //a1=8'd0
#560 a0=8'b10000000 ;a1=8'b00010000 ;a2=8'b00000000; //a2=8'd0
#610 a0=8'b10000000 ;a1=8'b00010000 ;a2=8'b00000011; //a2 error
#660 a0=8'b10000000 ;a1=8'b00010001 ;a2=8'b00000001; //a1 error
#710 a0=8'b10000001 ;a1=8'b00010000 ;a2=8'b00000001; //a0 error
#760 $finish;
end

initial $monitor ($time," a0=%d a1=%d a2=%d out=%d ",a0, a1, a2, out); 

// nwave
initial begin
	$fsdbDumpfile("median.fsdb");
	$fsdbDumpvars;
	$fsdbDumpMDA;
end

endmodule

